MOSFET Simulation
* this file edited to remove everything not in tt lib
.lib "./sky130_fd_pr/models/sky130.lib.spice" tt

X0 out input vdd vdd sky130_fd_pr__pfet_01v8 ad=3.06e+11p pd=2.26e+06u as=2.72e+11p ps=2.16e+06u w=680000u l=150000u
X1 out input VGND VGND sky130_fd_pr__nfet_01v8 ad=1.512e+11p pd=1.56e+06u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
C0 out vdd 0.06fF
C1 input vdd 0.07fF
C2 out input 0.02fF
C3 out VGND 0.13fF
C4 input VGND 0.25fF
C5 vdd VGND 0.55fF


* set gnd and power
Vgnd VGND 0 0
Vdd vdd VGND 1


* create pulse
Vin input VGND pulse(0 1 1p 10p 10p 1n 2n)
.tran 10p 2n 0

.control
run
set color0 = white
set color1 = black
plot input out
.endc

.end
